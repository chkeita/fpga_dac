module i2s_receiver_tb();
endmodule